module register_16_bit (
    input [15:0] D,     // 16-bit data input
    input clk,           // Clock input
    input rst,         // Asynchronous rst
    output [15:0] Q      // 16-bit data output
);

    // Create 16 D flip-flops for 16-bit register
    D_flip_flop DFF0 (.D(D[0]),   .clk(clk), .rst(rst), .Q(Q[0]));
    D_flip_flop DFF1 (.D(D[1]),   .clk(clk), .rst(rst), .Q(Q[1]));
    D_flip_flop DFF2 (.D(D[2]),   .clk(clk), .rst(rst), .Q(Q[2]));
    D_flip_flop DFF3 (.D(D[3]),   .clk(clk), .rst(rst), .Q(Q[3]));
    D_flip_flop DFF4 (.D(D[4]),   .clk(clk), .rst(rst), .Q(Q[4]));
    D_flip_flop DFF5 (.D(D[5]),   .clk(clk), .rst(rst), .Q(Q[5]));
    D_flip_flop DFF6 (.D(D[6]),   .clk(clk), .rst(rst), .Q(Q[6]));
    D_flip_flop DFF7 (.D(D[7]),   .clk(clk), .rst(rst), .Q(Q[7]));
    D_flip_flop DFF8 (.D(D[8]),   .clk(clk), .rst(rst), .Q(Q[8]));
    D_flip_flop DFF9 (.D(D[9]),   .clk(clk), .rst(rst), .Q(Q[9]));
    D_flip_flop DFF10 (.D(D[10]), .clk(clk), .rst(rst), .Q(Q[10]));
    D_flip_flop DFF11 (.D(D[11]), .clk(clk), .rst(rst), .Q(Q[11]));
    D_flip_flop DFF12 (.D(D[12]), .clk(clk), .rst(rst), .Q(Q[12]));
    D_flip_flop DFF13 (.D(D[13]), .clk(clk), .rst(rst), .Q(Q[13]));
    D_flip_flop DFF14 (.D(D[14]), .clk(clk), .rst(rst), .Q(Q[14]));
    D_flip_flop DFF15 (.D(D[15]), .clk(clk), .rst(rst), .Q(Q[15]));

endmodule
